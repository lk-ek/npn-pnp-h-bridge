
.model LED_3V D(IS=1e-13 RS=30 N=1.8 BV=5 CJO=0.2p IBV=10u)

.subckt LED_PAIR A B
R1 A N1 330
D1 N1 B LED_3V
R2 B N2 330
D2 N2 A LED_3V
.ends LED_PAIR

.subckt LED_ARRAY_14 A B
X1 A B LED_PAIR
X2 A B LED_PAIR
X3 A B LED_PAIR
X4 A B LED_PAIR
X5 A B LED_PAIR
X6 A B LED_PAIR
X7 A B LED_PAIR
X8 A B LED_PAIR
X9 A B LED_PAIR
X10 A B LED_PAIR
X11 A B LED_PAIR
X12 A B LED_PAIR
X13 A B LED_PAIR
X14 A B LED_PAIR
.ends LED_ARRAY_14

.subckt LED_ARRAY_28 A B
X1 A B LED_PAIR
X2 A B LED_PAIR
X3 A B LED_PAIR
X4 A B LED_PAIR
X5 A B LED_PAIR
X6 A B LED_PAIR
X7 A B LED_PAIR
X8 A B LED_PAIR
X9 A B LED_PAIR
X10 A B LED_PAIR
X11 A B LED_PAIR
X12 A B LED_PAIR
X13 A B LED_PAIR
X14 A B LED_PAIR
X15 A B LED_PAIR
X16 A B LED_PAIR
X17 A B LED_PAIR
X18 A B LED_PAIR
X19 A B LED_PAIR
X20 A B LED_PAIR
X21 A B LED_PAIR
X22 A B LED_PAIR
X23 A B LED_PAIR
X24 A B LED_PAIR
X25 A B LED_PAIR
X26 A B LED_PAIR
X27 A B LED_PAIR
X28 A B LED_PAIR
.ends LED_ARRAY_28

.subckt LED_ARRAY_42 A B
X1 A B LED_PAIR
X2 A B LED_PAIR
X3 A B LED_PAIR
X4 A B LED_PAIR
X5 A B LED_PAIR
X6 A B LED_PAIR
X7 A B LED_PAIR
X8 A B LED_PAIR
X9 A B LED_PAIR
X10 A B LED_PAIR
X11 A B LED_PAIR
X12 A B LED_PAIR
X13 A B LED_PAIR
X14 A B LED_PAIR
X15 A B LED_PAIR
X16 A B LED_PAIR
X17 A B LED_PAIR
X18 A B LED_PAIR
X19 A B LED_PAIR
X20 A B LED_PAIR
X21 A B LED_PAIR
X22 A B LED_PAIR
X23 A B LED_PAIR
X24 A B LED_PAIR
X25 A B LED_PAIR
X26 A B LED_PAIR
X27 A B LED_PAIR
X28 A B LED_PAIR
X29 A B LED_PAIR
X30 A B LED_PAIR
X31 A B LED_PAIR
X32 A B LED_PAIR
X33 A B LED_PAIR
X34 A B LED_PAIR
X35 A B LED_PAIR
X36 A B LED_PAIR
X37 A B LED_PAIR
X38 A B LED_PAIR
X39 A B LED_PAIR
X40 A B LED_PAIR
X41 A B LED_PAIR
X42 A B LED_PAIR
.ends LED_ARRAY_42

