
.model LED_3V D(IS=1e-13 RS=30 N=1.8 BV=5 CJO=0.2p IBV=10u)

.subckt LED_PAIR A B
R1 A N1 330
D1 N1 B LED_3V
R2 B N2 330
D2 N2 A LED_3V
.ends LED_PAIR

.subckt LED_ARRAY_2 A B
X1 A B LED_PAIR
X2 A B LED_PAIR
.ends LED_ARRAY_2

.subckt LED_ARRAY_4 A B
X1 A B LED_ARRAY_2
X2 A B LED_ARRAY_2
.ends LED_ARRAY_4

.subckt LED_ARRAY_8 A B
X1 A B LED_ARRAY_4
X2 A B LED_ARRAY_4
.ends LED_ARRAY_8

.subckt LED_ARRAY_14 A B
X1 A B LED_ARRAY_8
X2 A B LED_ARRAY_4
X3 A B LED_ARRAY_2
.ends LED_ARRAY_14

.subckt LED_ARRAY_16 A B
X1 A B LED_ARRAY_8
X2 A B LED_ARRAY_8
.ends LED_ARRAY_16

.subckt LED_ARRAY_28 A B
X1 A B LED_ARRAY_14
X2 A B LED_ARRAY_14
.ends LED_ARRAY_28

.subckt LED_ARRAY_32 A B
X1 A B LED_ARRAY_16
X2 A B LED_ARRAY_16
.ends LED_ARRAY_32

.subckt LED_ARRAY_42 A B
X1 A B LED_ARRAY_32
X2 A B LED_ARRAY_8
X3 A B LED_ARRAY_2
.ends LED_ARRAY_42

.subckt LED_ARRAY_64 A B
X1 A B LED_ARRAY_32
X2 A B LED_ARRAY_32
.ends LED_ARRAY_64

.subckt LED_ARRAY_84 A B
X1 A B LED_ARRAY_42
X2 A B LED_ARRAY_42
.ends LED_ARRAY_84

.subckt LED_ARRAY_128 A B
X1 A B LED_ARRAY_64
X2 A B LED_ARRAY_64
.ends LED_ARRAY_128

